module fifo_1 (input clock ,resetn,soft_reset,write_enb,read_enb,lfd_state,
        input [7:0]data_in , output reg[7:0]data_out, output full,empty);
integer count,i;
reg [4:0]wr_ptr,rd_ptr;
reg [8:0] mem [15:0];
reg lfd_reg;

always@(posedge clock)
	begin
		lfd_reg<=lfd_state;
	end

always@(posedge clock) //WRITE OPERATION
begin
	if(~resetn)
	begin
	for(i=0;i<16;i=i+1)
		mem[i]<=8'd0;
        end

	else if(soft_reset) //timeout condition,soft reset is generated by synchroniser
	       begin
		for(i=0;i<16;i=i+1)
			mem[i]<=8'd0;
	      end
	     
	
	     else 
                if(write_enb&&~full)
		{mem[wr_ptr[3:0]][8],mem[wr_ptr[3:0]][7:0]}<={lfd_reg,data_in};
	end
    

always@(posedge clock)
begin  
if(~resetn) data_out<=0;
else if(soft_reset) data_out<=8'dz;
else       
if(read_enb&&~empty)
		data_out<=mem[rd_ptr[3:0]][7:0];
end        
          
always@(posedge clock)
 begin 
 if(read_enb&&mem[rd_ptr[3:0]][8]&&~empty)
                count<=mem[rd_ptr[3:0]][7:2]+1'b1; //when ldf_state is 1, counter is loaded with payload lenght+1
	    else if(read_enb&&~mem[rd_ptr[3:0]][8] &&~empty)
		count<=count-1'b1;

		/*else if(count==0) data_out<=8'dz;

        end*/
end	

always@(posedge clock) //POINTER LOGIC
begin
	if(~resetn)
		wr_ptr<=0;
	if(soft_reset)
		wr_ptr<=0;
	else if(write_enb&&~full)
		wr_ptr<=wr_ptr+1'b1;
end
always @(posedge clock)
begin
	if(~resetn)
		rd_ptr<=0;
	if(soft_reset)
		rd_ptr<=0;
	else if(read_enb&&~empty)
		rd_ptr<=rd_ptr+1'b1;
end

assign empty=(rd_ptr==wr_ptr)?1'b1:1'b0;
assign full=((rd_ptr[4]!=wr_ptr[4])&&rd_ptr[3:0]==wr_ptr[3:0]);
endmodule
